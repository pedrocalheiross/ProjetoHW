module mux_DataSrc (
    input wire [31:0] data0, data1, data2, data3, data4, data5, data6, data7, data8,data9, data10, data11,
    input wire [1:0] AluSrcA, 
    output wire [31:0] out);


endmodule