module Controler(
    input wire clk,
    input wire reset,
    //...
);



endmodule